* Extracted by KLayout with SG13G2 LVS runset on : 29/04/2024 02:38

* cell sg13_lv_nmos
* pin sub!
.SUBCKT sg13_lv_nmos sub!
* device instance $1 r0 *1 3.765,-1.619 sg13_lv_nmos
M$1 \$6 \$12 \$1 sub! sg13_lv_nmos W=0.30000000000000004 L=0.3
* device instance $4 r0 *1 -0.059,-1.497 sg13_lv_nmos
M$4 \$3 \$8 \$5 sub! sg13_lv_nmos W=0.3 L=0.15
* device instance $6 r0 *1 0.023,0.275 sg13_lv_nmos
M$6 \$7 \$20 \$9 sub! sg13_lv_nmos W=0.15 L=0.13
* device instance $7 r0 *1 2.36,0.284 sg13_lv_nmos
M$7 \$10 \$24 \$11 sub! sg13_lv_nmos W=0.2 L=0.12999999999999998
* device instance $8 r0 *1 4.817,0.308 sg13_lv_nmos
M$8 \$16 \$26 \$17 sub! sg13_lv_nmos W=0.2 L=0.15
* device instance $9 r0 *1 0.02,2.078 sg13_lv_nmos
M$9 \$13 \$14 \$15 sub! sg13_lv_nmos W=0.6000000000000001 L=0.24999999999999997
* device instance $10 r0 *1 5.759,4.321 sg13_lv_nmos
M$10 \$27 \$29 \$19 sub! sg13_lv_nmos W=0.6 L=0.15
.ENDS sg13_lv_nmos
